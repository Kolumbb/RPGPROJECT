150 50
32
1
0 0 0 736 64 0 0 0 1 0 736 128 0 0 0 2 0 448 0 1 0 0 3 0 448 0 1 0 0 4 0 448 0 1 0 0 5 0 448 0 1 0 0 6 0 448 0 1 0 0 7 0 448 0 1 0 0 8 0 512 0 1 0 1 0 0 736 32 0 0 1 1 0 736 128 0 0 1 2 0 448 0 1 0 1 3 0 448 0 1 0 1 4 0 448 0 1 0 1 5 0 448 0 1 0 1 6 0 448 0 1 0 1 7 0 448 0 1 0 1 8 0 512 0 1 0 2 0 0 736 32 0 0 2 1 0 736 128 0 0 2 2 0 448 0 1 0 2 3 0 448 0 1 0 2 4 0 448 0 1 0 2 5 0 448 0 1 0 2 6 0 448 0 1 0 2 7 0 448 0 1 0 2 8 0 512 0 1 0 3 0 0 736 96 0 0 3 1 0 736 128 0 0 3 2 0 448 0 1 0 3 3 0 448 0 1 0 3 4 0 448 0 1 0 3 5 0 448 0 1 0 3 6 0 448 0 1 0 3 7 0 448 0 1 0 3 8 0 512 0 1 0 4 0 0 736 64 0 0 4 1 0 704 96 0 0 4 2 0 704 128 0 0 4 3 0 448 0 1 0 4 4 0 448 0 1 0 4 5 0 448 0 1 0 4 6 0 448 0 1 0 4 7 0 448 0 1 0 4 8 0 512 0 1 0 5 0 0 736 96 0 0 5 1 0 736 96 0 0 5 2 0 512 128 0 0 5 3 0 448 0 1 0 5 4 0 448 0 1 0 5 5 0 448 0 1 0 5 6 0 448 0 1 0 5 7 0 448 0 1 0 5 8 0 512 0 1 0 6 0 0 608 32 0 0 6 1 0 704 64 0 0 6 2 0 512 128 0 0 6 3 0 448 0 1 0 6 4 0 448 0 1 0 6 5 0 448 0 1 0 6 6 0 448 0 1 0 6 7 0 448 0 1 0 6 8 0 512 0 1 0 7 0 0 736 0 0 0 7 1 0 704 64 0 0 7 2 0 512 128 0 0 7 3 0 448 0 1 0 7 4 0 448 0 1 0 7 5 0 448 0 1 0 7 6 0 448 0 1 0 7 7 0 448 0 1 0 7 8 0 512 0 1 0 7 9 0 32 64 0 0 7 10 0 32 64 0 0 7 11 0 736 64 0 0 7 12 0 736 64 0 0 7 13 0 736 64 0 0 7 14 0 736 64 0 0 7 15 0 288 32 0 0 7 16 0 288 32 0 0 7 17 0 288 32 0 0 7 18 0 736 64 0 0 7 19 0 288 32 0 0 7 20 0 288 32 0 0 7 21 0 736 64 0 0 7 22 0 736 64 0 0 7 23 0 736 64 0 0 7 24 0 736 64 0 0 7 25 0 736 64 0 0 7 26 0 736 64 0 0 7 27 0 736 64 0 0 7 28 0 736 64 0 0 7 29 0 736 64 0 0 7 30 0 736 64 0 0 7 31 0 736 64 0 0 7 32 0 736 64 0 0 7 33 0 736 64 0 0 8 0 0 736 0 0 0 8 1 0 736 96 0 0 8 2 0 512 128 0 0 8 3 0 448 0 1 0 8 4 0 448 0 1 0 8 5 0 448 0 1 0 8 6 0 448 0 1 0 8 7 0 480 0 1 0 8 8 0 480 32 1 0 8 9 0 736 64 0 0 8 10 0 736 64 0 0 8 11 0 736 64 0 0 8 12 0 736 64 0 0 8 13 0 736 64 0 0 8 14 0 736 64 0 0 8 15 0 32 64 0 0 8 16 0 32 64 0 0 8 17 0 736 64 0 0 8 18 0 736 64 0 0 8 19 0 288 32 0 0 8 20 0 736 64 0 0 8 21 0 736 64 0 0 8 22 0 32 64 0 0 8 23 0 32 64 0 0 8 24 0 736 64 0 0 8 25 0 32 64 0 0 8 26 0 736 64 0 0 8 27 0 736 64 0 0 8 28 0 736 64 0 0 8 29 0 736 64 0 0 8 30 0 736 64 0 0 8 31 0 736 64 0 0 8 32 0 736 64 0 0 8 33 0 736 64 0 0 9 0 0 736 0 0 0 9 1 0 704 64 0 0 9 2 0 512 128 0 0 9 3 0 448 0 1 0 9 4 0 448 0 1 0 9 5 0 448 0 1 0 9 6 0 448 0 1 0 9 7 0 512 0 1 0 9 8 0 320 64 0 0 9 9 0 736 64 0 0 9 10 0 32 64 0 0 9 11 0 736 64 0 0 9 12 0 736 64 0 0 9 13 0 736 64 0 0 9 14 0 736 64 0 0 9 15 0 288 32 0 0 9 16 0 736 64 0 0 9 17 0 736 64 0 0 9 18 0 736 64 0 0 9 19 0 32 64 0 0 9 20 0 32 64 0 0 9 21 0 736 64 0 0 9 22 0 736 64 0 0 9 23 0 32 64 0 0 9 24 0 32 64 0 0 9 25 0 736 64 0 0 9 26 0 736 64 0 0 9 27 0 736 64 0 0 9 28 0 736 64 0 0 9 29 0 736 64 0 0 9 30 0 736 64 0 0 9 31 0 736 64 0 0 9 32 0 736 64 0 0 9 33 0 736 64 0 0 10 0 0 640 32 0 0 10 1 0 704 64 0 0 10 2 0 512 128 0 0 10 3 0 448 0 1 0 10 4 0 448 0 1 0 10 5 0 448 0 1 0 10 6 0 448 0 1 0 10 7 0 512 0 1 0 10 8 0 736 64 0 0 10 9 0 736 64 0 0 10 10 0 736 64 0 0 10 11 0 736 64 0 0 10 12 0 736 64 0 0 10 13 0 736 64 0 0 10 14 0 32 64 0 0 10 15 0 288 32 0 0 10 16 0 736 64 0 0 10 17 0 32 64 0 0 10 18 0 32 64 0 0 10 19 0 288 32 0 0 10 20 0 736 64 0 0 10 21 0 736 64 0 0 10 22 0 736 64 0 0 10 23 0 736 64 0 0 10 24 0 736 64 0 0 10 25 0 736 64 0 0 10 26 0 32 64 0 0 10 27 0 736 64 0 0 10 28 0 736 64 0 0 10 29 0 736 64 0 0 10 30 0 736 64 0 0 10 31 0 736 64 0 0 10 32 0 736 64 0 0 10 33 0 736 64 0 0 11 0 0 704 64 0 0 11 1 0 736 96 0 0 11 2 0 512 128 0 0 11 3 0 448 0 1 0 11 4 0 448 0 1 0 11 5 0 448 0 1 0 11 6 0 448 0 1 0 11 7 0 512 0 1 0 11 8 0 736 64 0 0 11 9 0 736 64 0 0 11 10 0 256 64 0 0 11 11 0 256 64 0 0 11 12 0 736 64 0 0 11 13 0 736 64 0 0 11 14 0 736 64 0 0 11 15 0 288 32 0 0 11 16 0 768 64 0 0 11 17 0 32 64 0 0 11 18 0 288 32 0 0 11 19 0 288 32 0 0 11 20 0 64 32 0 0 11 21 0 768 64 0 0 11 22 0 736 64 0 0 11 23 0 32 64 0 0 11 24 0 32 64 0 0 11 25 0 736 64 0 0 11 26 0 32 64 0 0 11 27 0 736 64 0 0 11 28 0 736 64 0 0 11 29 0 736 64 0 0 11 30 0 736 64 0 0 11 31 0 736 64 0 0 11 32 0 736 64 0 0 11 33 0 736 64 0 0 12 0 0 800 64 0 0 12 1 0 800 64 0 0 12 2 0 768 128 0 0 12 3 0 448 0 1 0 12 4 0 448 0 1 0 12 5 0 448 0 1 0 12 6 0 448 0 1 0 12 7 0 512 0 1 0 12 8 0 736 64 0 0 12 9 0 736 64 0 0 12 10 0 736 64 0 0 12 11 0 736 64 0 0 12 12 0 288 32 0 0 12 13 0 288 32 0 0 12 14 0 320 64 0 0 12 15 0 320 64 0 0 12 16 0 736 64 0 0 12 17 0 736 64 0 0 12 18 0 288 32 0 0 12 19 0 736 64 0 0 12 20 0 736 64 0 0 12 21 0 736 64 0 0 12 22 0 736 64 0 0 12 23 0 64 32 0 0 12 24 0 32 64 0 0 12 25 0 736 64 0 0 12 26 0 32 64 0 0 12 27 0 736 64 0 0 12 28 0 32 64 0 0 12 29 0 32 64 0 0 12 30 0 32 64 0 0 12 31 0 736 64 0 0 12 32 0 736 64 0 0 12 33 0 736 64 0 0 13 0 0 448 0 1 0 13 1 0 448 0 1 0 13 2 0 448 0 1 0 13 3 0 448 0 1 0 13 4 0 448 0 1 0 13 5 0 448 0 1 0 13 6 0 448 0 1 0 13 7 0 512 0 1 0 13 8 0 736 64 0 0 13 9 0 96 64 0 0 13 10 0 32 64 0 0 13 11 0 96 64 0 0 13 12 0 288 32 0 0 13 13 0 96 64 0 0 13 14 0 96 64 0 0 13 15 0 320 64 0 0 13 16 0 736 64 0 0 13 17 0 96 64 0 0 13 18 0 288 32 0 0 13 19 0 288 32 0 0 13 20 0 736 64 0 0 13 21 0 480 64 0 0 13 22 0 736 64 0 0 13 23 0 64 32 0 0 13 24 0 32 64 0 0 13 25 0 736 64 0 0 13 26 0 32 64 0 0 13 27 0 32 64 0 0 13 28 0 32 64 0 0 13 29 0 32 64 0 0 13 30 0 736 64 0 0 13 31 0 32 64 0 0 13 32 0 736 64 0 0 13 33 0 736 64 0 0 14 0 0 448 0 1 0 14 1 0 448 0 1 0 14 2 0 448 0 1 0 14 3 0 448 0 1 0 14 4 0 448 0 1 0 14 5 0 448 0 1 0 14 6 0 480 0 1 0 14 7 0 480 32 1 0 14 8 0 256 64 0 0 14 9 0 96 64 0 0 14 10 0 256 64 0 0 14 11 0 736 64 0 0 14 12 0 288 32 0 0 14 13 0 320 64 0 0 14 14 0 736 64 0 0 14 15 0 736 64 0 0 14 16 0 736 64 0 0 14 17 0 736 64 0 0 14 18 0 736 64 0 0 14 19 0 96 64 0 0 14 20 0 288 32 0 0 14 21 0 480 64 0 0 14 22 0 480 64 0 0 14 23 0 64 32 0 0 14 24 0 736 64 0 0 14 25 0 736 64 0 0 14 26 0 32 64 0 0 14 27 0 32 64 0 0 14 28 0 736 64 0 0 14 29 0 32 64 0 0 14 30 0 32 64 0 0 14 31 0 32 64 0 0 14 32 0 32 64 0 0 14 33 0 736 64 0 0 15 0 0 448 0 1 0 15 1 0 448 0 1 0 15 2 0 448 0 1 0 15 3 0 448 0 1 0 15 4 0 448 0 1 0 15 5 0 448 0 1 0 15 6 0 512 0 1 0 15 7 0 256 64 0 0 15 8 0 736 64 0 0 15 9 0 96 64 0 0 15 10 0 736 64 0 0 15 11 0 96 96 1 1 15 12 0 736 64 0 0 15 13 0 736 64 0 0 15 14 0 736 64 0 0 15 15 0 768 64 0 0 15 16 0 320 64 0 0 15 17 0 64 32 0 0 15 18 0 736 64 0 0 15 19 0 288 32 0 0 15 20 0 736 64 0 0 15 21 0 736 64 0 0 15 22 0 480 64 0 0 15 23 0 64 32 0 0 15 24 0 736 64 0 0 15 25 0 32 64 0 0 15 26 0 32 64 0 0 15 27 0 32 64 0 0 15 28 0 32 64 0 0 15 29 0 32 64 0 0 15 30 0 736 64 0 0 15 31 0 32 64 0 0 15 32 0 32 64 0 0 15 33 0 736 64 0 0 16 0 0 448 64 1 0 16 1 0 448 64 1 0 16 2 0 448 64 1 0 16 3 0 448 64 1 0 16 4 0 448 64 1 0 16 5 0 448 64 1 0 16 6 0 480 32 1 0 16 7 0 256 64 0 0 16 8 0 736 64 0 0 16 9 0 96 64 0 0 16 10 0 768 64 0 0 16 11 0 736 64 0 0 16 12 0 288 32 0 0 16 13 0 736 64 0 0 16 14 0 288 96 0 0 16 15 0 736 64 0 0 16 16 0 320 64 0 0 16 17 0 288 96 0 0 16 18 0 288 96 0 0 16 19 0 288 96 0 0 16 20 0 736 64 0 0 16 21 0 288 96 0 0 16 22 0 480 64 0 0 16 23 0 64 32 0 0 16 24 0 736 64 0 0 16 25 0 736 64 0 0 16 26 0 736 64 0 0 16 27 0 32 64 0 0 16 28 0 32 64 0 0 16 29 0 32 64 0 0 16 30 0 736 64 0 0 16 31 0 32 64 0 0 16 32 0 736 64 0 0 16 33 0 736 64 0 0 17 0 0 736 64 0 0 17 1 0 480 64 0 0 17 2 0 736 64 0 0 17 3 0 256 64 0 0 17 4 0 736 64 0 0 17 5 0 736 64 0 0 17 6 0 736 64 0 0 17 7 0 256 64 0 0 17 8 0 736 64 0 0 17 9 0 96 64 0 0 17 10 0 64 32 0 0 17 11 0 64 32 0 0 17 12 0 288 32 0 0 17 13 0 320 64 0 0 17 14 0 320 64 0 0 17 15 0 320 64 0 0 17 16 0 320 64 0 0 17 17 0 480 64 0 0 17 18 0 480 64 0 0 17 19 0 480 64 0 0 17 20 0 480 64 0 0 17 21 0 768 64 0 0 17 22 0 288 96 0 0 17 23 0 480 64 0 0 17 24 0 64 32 0 0 17 25 0 736 64 0 0 17 26 0 64 32 0 0 17 27 0 736 64 0 0 17 28 0 736 64 0 0 17 29 0 64 32 0 0 17 30 0 64 32 0 0 17 31 0 32 64 0 0 17 32 0 32 64 0 0 17 33 0 736 64 0 0 18 0 0 480 64 0 0 18 1 0 480 64 0 0 18 2 0 736 64 0 0 18 3 0 480 64 0 0 18 4 0 704 64 0 0 18 5 0 736 64 0 0 18 6 0 736 64 0 0 18 7 0 256 64 0 0 18 8 0 736 64 0 0 18 9 0 288 32 0 0 18 10 0 288 32 0 0 18 11 0 288 32 0 0 18 12 0 320 64 0 0 18 13 0 320 64 0 0 18 14 0 736 64 0 0 18 15 0 480 64 0 0 18 16 0 736 64 0 0 18 17 0 320 64 0 0 18 18 0 96 64 0 0 18 19 0 288 96 0 0 18 20 0 96 64 0 0 18 21 0 288 96 0 0 18 22 0 736 64 0 0 18 23 0 480 64 0 0 18 24 0 736 64 0 0 18 25 0 736 64 0 0 18 26 0 64 32 0 0 18 27 0 736 64 0 0 18 28 0 64 32 0 0 18 29 0 736 64 0 0 18 30 0 736 64 0 0 18 31 0 64 32 0 0 18 32 0 736 64 0 0 18 33 0 736 64 0 0 19 0 0 288 32 0 0 19 1 0 64 32 0 0 19 2 0 64 32 0 0 19 3 0 736 64 0 0 19 4 0 704 64 0 0 19 5 0 736 64 0 0 19 6 0 736 64 0 0 19 7 0 736 64 0 0 19 8 0 736 64 0 0 19 9 0 288 32 0 0 19 10 0 736 64 0 0 19 11 0 736 64 0 0 19 12 0 320 64 0 0 19 13 0 736 64 0 0 19 14 0 288 96 0 0 19 15 0 96 64 0 0 19 16 0 736 64 0 0 19 17 0 320 64 0 0 19 18 0 768 64 0 0 19 19 0 288 96 0 0 19 20 0 288 96 0 0 19 21 0 480 64 0 0 19 22 0 480 64 0 0 19 23 0 288 96 0 0 19 24 0 288 96 0 0 19 25 0 736 64 0 0 19 26 0 64 32 0 0 19 27 0 736 64 0 0 19 28 0 64 32 0 0 19 29 0 736 64 0 0 19 30 0 32 64 0 0 19 31 0 64 32 0 0 19 32 0 32 64 0 0 19 33 0 736 64 0 0 20 0 0 64 32 0 0 20 1 0 736 64 0 0 20 2 0 64 32 0 0 20 3 0 480 64 0 0 20 4 0 736 64 0 0 20 5 0 736 64 0 0 20 6 0 736 64 0 0 20 7 0 736 64 0 0 20 8 0 768 64 0 0 20 9 0 288 32 0 0 20 10 0 288 32 0 0 20 11 0 288 32 0 0 20 12 0 320 64 0 0 20 13 0 288 32 0 0 20 14 0 288 96 0 0 20 15 0 768 64 0 0 20 16 0 288 96 0 0 20 17 0 736 64 0 0 20 18 0 320 64 0 0 20 19 0 480 64 0 0 20 20 0 288 96 0 0 20 21 0 320 64 0 0 20 22 0 320 64 0 0 20 23 0 736 64 0 0 20 24 0 288 96 0 0 20 25 0 736 64 0 0 20 26 0 736 64 0 0 20 27 0 64 32 0 0 20 28 0 64 32 0 0 20 29 0 736 64 0 0 20 30 0 32 64 0 0 20 31 0 64 32 0 0 20 32 0 736 64 0 0 20 33 0 736 64 0 0 21 0 0 736 64 0 0 21 1 0 736 64 0 0 21 2 0 736 64 0 0 21 3 0 736 64 0 0 21 4 0 736 64 0 0 21 5 0 736 64 0 0 21 6 0 736 64 0 0 21 7 0 736 64 0 0 21 8 0 736 64 0 0 21 9 0 320 64 0 0 21 10 0 736 64 0 0 21 11 0 736 64 0 0 21 12 0 768 64 0 0 21 13 0 288 32 0 0 21 14 0 288 96 0 0 21 15 0 96 64 0 0 21 16 0 480 64 0 0 21 17 0 320 64 0 0 21 18 0 320 64 0 0 21 19 0 736 64 0 0 21 20 0 480 64 0 0 21 21 0 480 64 0 0 21 22 0 480 64 0 0 21 23 0 480 64 0 0 21 24 0 288 96 0 0 21 25 0 736 64 0 0 21 26 0 736 64 0 0 21 27 0 64 32 0 0 21 28 0 64 32 0 0 21 29 0 64 32 0 0 21 30 0 64 32 0 0 21 31 0 736 64 0 0 21 32 0 736 64 0 0 21 33 0 736 64 0 0 22 0 0 480 64 0 0 22 1 0 736 64 0 0 22 2 0 480 64 0 0 22 3 0 480 64 0 0 22 4 0 736 64 0 0 22 5 0 736 64 0 0 22 6 0 736 64 0 0 22 7 0 256 64 0 0 22 8 0 256 64 0 0 22 9 0 256 64 0 0 22 10 0 256 64 0 0 22 11 0 256 64 0 0 22 12 0 256 64 0 0 22 13 0 288 32 0 0 22 14 0 288 32 0 0 22 15 0 288 96 0 0 22 16 0 480 64 0 0 22 17 0 288 96 0 0 22 18 0 288 32 0 0 22 19 0 288 32 0 0 22 20 0 736 64 0 0 22 21 0 768 64 0 0 22 22 0 96 64 0 0 22 23 0 480 64 0 0 22 24 0 96 64 0 0 22 25 0 64 32 0 0 22 26 0 64 32 0 0 22 27 0 64 32 0 0 22 28 0 64 32 0 0 22 29 0 64 32 0 0 22 30 0 64 32 0 0 22 31 0 736 64 0 0 22 32 0 736 64 0 0 22 33 0 736 64 0 0 23 0 0 64 32 0 0 23 1 0 736 64 0 0 23 2 0 64 32 0 0 23 3 0 288 32 0 0 23 4 0 480 64 0 0 23 5 0 736 64 0 0 23 6 0 736 64 0 0 23 7 0 736 64 0 0 23 8 0 736 64 0 0 23 9 0 96 64 0 0 23 10 0 480 64 0 0 23 11 0 736 64 0 0 23 12 0 320 64 0 0 23 13 0 480 64 0 0 23 14 0 768 64 0 0 23 15 0 96 64 0 0 23 16 0 288 32 0 0 23 17 0 736 64 0 0 23 18 0 288 32 0 0 23 19 0 736 64 0 0 23 20 0 320 64 0 0 23 21 0 96 64 0 0 23 22 0 320 64 0 0 23 23 0 736 64 0 0 23 24 0 288 96 0 0 23 25 0 64 32 0 0 23 26 0 736 64 0 0 23 27 0 64 32 0 0 23 28 0 64 32 0 0 23 29 0 736 64 0 0 23 30 0 64 32 0 0 23 31 0 64 32 0 0 23 32 0 736 64 0 0 23 33 0 736 64 0 0 24 0 0 288 32 0 0 24 1 0 288 32 0 0 24 2 0 64 32 0 0 24 3 0 64 32 0 0 24 4 0 736 64 0 0 24 5 0 736 64 0 0 24 6 0 768 64 0 0 24 7 0 768 64 0 0 24 8 0 768 64 0 0 24 9 0 768 64 0 0 24 10 0 736 64 0 0 24 11 0 736 64 0 0 24 12 0 480 64 0 0 24 13 0 736 64 0 0 24 14 0 288 96 0 0 24 15 0 480 64 0 0 24 16 0 288 32 0 0 24 17 0 736 64 0 0 24 18 0 736 64 0 0 24 19 0 320 64 0 0 24 20 0 320 64 0 0 24 21 0 96 64 0 0 24 22 0 320 64 0 0 24 23 0 736 64 0 0 24 24 0 64 32 0 0 24 25 0 736 64 0 0 24 26 0 96 64 0 0 24 27 0 736 64 0 0 24 28 0 736 64 0 0 24 29 0 736 64 0 0 24 30 0 736 64 0 0 24 31 0 64 32 0 0 24 32 0 736 64 0 0 24 33 0 736 64 0 0 25 0 0 288 32 0 0 25 1 0 288 32 0 0 25 2 0 64 32 0 0 25 3 0 64 32 0 0 25 4 0 704 64 0 0 25 5 0 736 64 0 0 25 6 0 736 64 0 0 25 7 0 736 64 0 0 25 8 0 736 64 0 0 25 9 0 736 64 0 0 25 10 0 512 96 0 0 25 11 0 736 64 0 0 25 12 0 288 32 0 0 25 13 0 736 64 0 0 25 14 0 736 64 0 0 25 15 0 480 64 0 0 25 16 0 736 64 0 0 25 17 0 736 64 0 0 25 18 0 320 64 0 0 25 19 0 320 64 0 0 25 20 0 768 64 0 0 25 21 0 544 64 0 0 25 22 0 320 64 0 0 25 23 0 736 64 0 0 25 24 0 288 96 0 0 25 25 0 736 64 0 0 25 26 0 96 64 0 0 25 27 0 96 64 0 0 25 28 0 64 32 0 0 25 29 0 736 64 0 0 25 30 0 736 64 0 0 25 31 0 64 32 0 0 25 32 0 736 64 0 0 25 33 0 736 64 0 0 26 0 0 736 64 0 0 26 1 0 288 32 0 0 26 2 0 736 64 0 0 26 3 0 288 32 0 0 26 4 0 480 64 0 0 26 5 0 736 64 0 0 26 6 0 736 64 0 0 26 7 0 736 64 0 0 26 8 0 736 64 0 0 26 9 0 512 96 0 0 26 10 0 736 64 0 0 26 11 0 736 64 0 0 26 12 0 288 32 0 0 26 13 0 512 96 0 0 26 14 0 736 64 0 0 26 15 0 736 64 0 0 26 16 0 768 64 0 0 26 17 0 768 64 0 0 26 18 0 544 64 0 0 26 19 0 736 64 0 0 26 20 0 736 64 0 0 26 21 0 736 64 0 0 26 22 0 320 64 0 0 26 23 0 736 64 0 0 26 24 0 288 96 0 0 26 25 0 736 64 0 0 26 26 0 736 64 0 0 26 27 0 96 64 0 0 26 28 0 736 64 0 0 26 29 0 736 64 0 0 26 30 0 64 32 0 0 26 31 0 64 32 0 0 26 32 0 736 64 0 0 26 33 0 736 64 0 0 27 0 0 736 64 0 0 27 1 0 480 64 0 0 27 2 0 64 32 0 0 27 3 0 736 64 0 0 27 4 0 704 64 0 0 27 5 0 736 64 0 0 27 6 0 736 64 0 0 27 7 0 736 64 0 0 27 8 0 736 64 0 0 27 9 0 512 96 0 0 27 10 0 320 64 0 0 27 11 0 736 64 0 0 27 12 0 288 32 0 0 27 13 0 512 96 0 0 27 14 0 512 96 0 0 27 15 0 768 64 0 0 27 16 0 736 64 0 0 27 17 0 736 64 0 0 27 18 0 320 64 0 0 27 19 0 288 32 0 0 27 20 0 288 32 0 0 27 21 0 544 64 0 0 27 22 0 288 32 0 0 27 23 0 288 32 0 0 27 24 0 288 96 0 0 27 25 0 736 64 0 0 27 26 0 736 64 0 0 27 27 0 736 64 0 0 27 28 0 96 64 0 0 27 29 0 96 64 0 0 27 30 0 736 64 0 0 27 31 0 736 64 0 0 27 32 0 736 64 0 0 27 33 0 736 64 0 0 28 0 0 704 64 0 0 28 1 0 480 64 0 0 28 2 0 64 32 0 0 28 3 0 64 32 0 0 28 4 0 704 64 0 0 28 5 0 736 64 0 0 28 6 0 736 64 0 0 28 7 0 736 64 0 0 28 8 0 736 64 0 0 28 9 0 736 64 0 0 28 10 0 736 64 0 0 28 11 0 736 64 0 0 28 12 0 736 64 0 0 28 13 0 736 64 0 0 28 14 0 512 96 0 0 28 15 0 512 96 0 0 28 16 0 768 64 0 0 28 17 0 768 64 0 0 28 18 0 768 64 0 0 28 19 0 768 64 0 0 28 20 0 288 32 0 0 28 21 0 736 64 0 0 28 22 0 736 64 0 0 28 23 0 320 64 0 0 28 24 0 288 96 0 0 28 25 0 736 64 0 0 28 26 0 736 64 0 0 28 27 0 96 64 0 0 28 28 0 96 64 0 0 28 29 0 736 64 0 0 28 30 0 736 64 0 0 28 31 0 736 64 0 0 28 32 0 736 64 0 0 28 33 0 736 64 0 0 29 0 0 288 32 0 0 29 1 0 736 64 0 0 29 2 0 704 64 0 0 29 3 0 64 32 0 0 29 4 0 64 32 0 0 29 5 0 736 64 0 0 29 6 0 736 64 0 0 29 7 0 736 64 0 0 29 8 0 320 64 0 0 29 9 0 320 64 0 0 29 10 0 736 64 0 0 29 11 0 512 96 0 0 29 12 0 736 64 0 0 29 13 0 288 96 0 0 29 14 0 736 64 0 0 29 15 0 736 64 0 0 29 16 0 512 96 0 0 29 17 0 736 64 0 0 29 18 0 736 64 0 0 29 19 0 320 64 0 0 29 20 0 320 64 0 0 29 21 0 64 32 0 0 29 22 0 320 64 0 0 29 23 0 320 64 0 0 29 24 0 288 96 0 0 29 25 0 64 32 0 0 29 26 0 736 64 0 0 29 27 0 96 64 0 0 29 28 0 64 32 0 0 29 29 0 736 64 0 0 29 30 0 736 64 0 0 29 31 0 736 64 0 0 29 32 0 736 64 0 0 29 33 0 736 64 0 0 30 0 0 704 64 0 0 30 1 0 64 32 0 0 30 2 0 704 64 0 0 30 3 0 64 32 0 0 30 4 0 704 64 0 0 30 5 0 736 64 0 0 30 6 0 736 64 0 0 30 7 0 288 32 0 0 30 8 0 320 64 0 0 30 9 0 736 64 0 0 30 10 0 512 352 0 1 30 11 0 320 64 0 0 30 12 0 320 64 0 0 30 13 0 288 32 0 0 30 14 0 288 32 0 0 30 15 0 288 32 0 0 30 16 0 320 64 0 0 30 17 0 512 96 0 0 30 18 0 768 64 0 0 30 19 0 512 96 0 0 30 20 0 512 96 0 0 30 21 0 736 64 0 0 30 22 0 512 96 0 0 30 23 0 736 64 0 0 30 24 0 288 96 0 0 30 25 0 736 64 0 0 30 26 0 96 64 0 0 30 27 0 96 64 0 0 30 28 0 64 32 0 0 30 29 0 736 64 0 0 30 30 0 736 64 0 0 30 31 0 736 64 0 0 30 32 0 736 64 0 0 30 33 0 736 64 0 0 31 0 0 704 64 0 0 31 1 0 288 32 0 0 31 2 0 64 32 0 0 31 3 0 288 32 0 0 31 4 0 704 64 0 0 31 5 0 736 64 0 0 31 6 0 736 64 0 0 31 7 0 736 64 0 0 31 8 0 736 64 0 0 31 9 0 288 32 0 0 31 10 0 736 64 0 0 31 11 0 512 96 0 0 31 12 0 736 64 0 0 31 13 0 736 64 0 0 31 14 0 736 64 0 0 31 15 0 736 64 0 0 31 16 0 736 64 0 0 31 17 0 768 64 0 0 31 18 0 288 96 0 0 31 19 0 736 64 0 0 31 20 0 288 96 0 0 31 21 0 736 64 0 0 31 22 0 64 32 0 0 31 23 0 64 32 0 0 31 24 0 288 96 0 0 31 25 0 96 64 0 0 31 26 0 96 64 0 0 31 27 0 736 64 0 0 31 28 0 736 64 0 0 31 29 0 736 64 0 0 31 30 0 736 64 0 0 31 31 0 736 64 0 0 31 32 0 736 64 0 0 31 33 0 736 64 0 0 32 0 0 288 32 0 0 32 1 0 288 32 0 0 32 2 0 704 64 0 0 32 3 0 736 64 0 0 32 4 0 64 32 0 0 32 5 0 288 32 0 0 32 6 0 736 64 0 0 32 7 0 736 64 0 0 32 8 0 736 64 0 0 32 9 0 736 64 0 0 32 10 0 736 64 0 0 32 11 0 736 64 0 0 32 12 0 736 64 0 0 32 13 0 512 96 0 0 32 14 0 512 96 0 0 32 15 0 736 64 0 0 32 16 0 320 64 0 0 32 17 0 320 64 0 0 32 18 0 736 64 0 0 32 19 0 736 64 0 0 32 20 0 320 64 0 0 32 21 0 320 64 0 0 32 22 0 736 64 0 0 32 23 0 288 96 0 0 32 24 0 96 64 0 0 32 25 0 96 64 0 0 32 26 0 736 64 0 0 32 27 0 736 64 0 0 32 28 0 736 64 0 0 32 29 0 736 64 0 0 32 30 0 736 64 0 0 32 31 0 736 64 0 0 32 32 0 736 64 0 0 32 33 0 736 64 0 0 33 0 0 704 64 0 0 33 1 0 480 64 0 0 33 2 0 736 64 0 0 33 3 0 736 64 0 0 33 4 0 736 64 0 0 33 5 0 736 64 0 0 33 6 0 288 32 0 0 33 7 0 736 64 0 0 33 8 0 736 64 0 0 33 9 0 736 64 0 0 33 10 0 736 64 0 0 33 11 0 736 64 0 0 33 12 0 320 64 0 0 33 13 0 736 64 0 0 33 14 0 736 64 0 0 33 15 0 736 64 0 0 33 16 0 320 64 0 0 33 17 0 736 64 0 0 33 18 0 320 64 0 0 33 19 0 736 64 0 0 33 20 0 288 32 0 0 33 21 0 320 64 0 0 33 22 0 736 64 0 0 33 23 0 64 32 0 0 33 24 0 736 64 0 0 33 25 0 736 64 0 0 33 26 0 736 64 0 0 33 27 0 736 64 0 0 33 28 0 736 64 0 0 33 29 0 736 64 0 0 33 30 0 736 64 0 0 33 31 0 736 64 0 0 33 32 0 736 64 0 0 33 33 0 736 64 0 0 34 0 0 704 64 0 0 34 1 0 288 32 0 0 34 2 0 736 64 0 0 34 3 0 736 64 0 0 34 4 0 64 32 0 0 34 5 0 736 64 0 0 34 6 0 736 64 0 0 34 7 0 736 64 0 0 34 8 0 736 64 0 0 34 9 0 288 32 0 0 34 10 0 736 64 0 0 34 11 0 96 64 0 0 34 12 0 320 64 0 0 34 13 0 96 64 0 0 34 14 0 736 64 0 0 34 15 0 96 64 0 0 34 16 0 320 64 0 0 34 17 0 736 64 0 0 34 18 0 736 64 0 0 34 19 0 768 64 0 0 34 20 0 736 64 0 0 34 21 0 736 64 0 0 34 22 0 736 64 0 0 34 23 0 736 64 0 0 34 24 0 736 64 0 0 34 25 0 736 64 0 0 34 26 0 736 64 0 0 34 27 0 736 64 0 0 34 28 0 736 64 0 0 34 29 0 736 64 0 0 34 30 0 736 64 0 0 34 31 0 736 64 0 0 34 32 0 736 64 0 0 34 33 0 736 64 0 0 35 0 0 288 32 0 0 35 1 0 64 32 0 0 35 2 0 288 32 0 0 35 3 0 704 64 0 0 35 4 0 480 64 0 0 35 5 0 736 64 0 0 35 6 0 736 64 0 0 35 7 0 736 64 0 0 35 8 0 736 64 0 0 35 9 0 736 64 0 0 35 10 0 736 64 0 0 35 11 0 736 64 0 0 35 12 0 736 64 0 0 35 13 0 736 64 0 0 35 14 0 736 64 0 0 35 15 0 320 64 0 0 35 16 0 288 32 0 0 35 17 0 736 64 0 0 35 18 0 736 64 0 0 35 19 0 736 64 0 0 35 20 0 736 64 0 0 35 21 0 736 64 0 0 35 22 0 736 64 0 0 35 23 0 736 64 0 0 35 24 0 736 64 0 0 35 25 0 736 64 0 0 35 26 0 736 64 0 0 35 27 0 736 64 0 0 35 28 0 736 64 0 0 35 29 0 736 64 0 0 35 30 0 736 64 0 0 35 31 0 736 64 0 0 35 32 0 736 64 0 0 35 33 0 736 64 0 0 36 0 0 704 64 0 0 36 1 0 64 32 0 0 36 2 0 288 32 0 0 36 3 0 64 32 0 0 36 4 0 480 64 0 0 36 5 0 736 64 0 0 36 6 0 736 64 0 0 36 7 0 736 64 0 0 36 8 0 736 64 0 0 36 9 0 736 64 0 0 36 10 0 736 64 0 0 36 11 0 736 64 0 0 36 12 0 320 64 0 0 36 13 0 320 64 0 0 36 14 0 736 64 0 0 36 15 0 736 64 0 0 36 16 0 736 64 0 0 36 17 0 736 64 0 0 36 18 0 736 64 0 0 36 19 0 736 64 0 0 36 20 0 736 64 0 0 36 21 0 736 64 0 0 36 22 0 736 64 0 0 36 23 0 736 64 0 0 36 24 0 736 64 0 0 36 25 0 736 64 0 0 36 26 0 736 64 0 0 36 27 0 736 64 0 0 36 28 0 736 64 0 0 36 29 0 736 64 0 0 36 30 0 736 64 0 0 36 31 0 736 64 0 0 36 32 0 736 64 0 0 36 33 0 736 64 0 0 37 0 0 704 64 0 0 37 1 0 64 32 0 0 37 2 0 288 32 0 0 37 3 0 64 32 0 0 37 4 0 64 32 0 0 37 5 0 736 64 0 0 37 6 0 736 64 0 0 37 7 0 736 64 0 0 37 8 0 736 64 0 0 37 9 0 736 64 0 0 37 10 0 736 64 0 0 37 11 0 736 64 0 0 37 12 0 736 64 0 0 37 13 0 736 64 0 0 37 14 0 736 64 0 0 37 15 0 736 64 0 0 37 16 0 736 64 0 0 37 17 0 736 64 0 0 37 18 0 736 64 0 0 37 19 0 736 64 0 0 37 20 0 736 64 0 0 37 21 0 736 64 0 0 37 22 0 736 64 0 0 37 23 0 736 64 0 0 37 24 0 736 64 0 0 37 25 0 736 64 0 0 37 26 0 736 64 0 0 37 27 0 736 64 0 0 37 28 0 736 64 0 0 37 29 0 736 64 0 0 37 30 0 736 64 0 0 37 31 0 736 64 0 0 37 32 0 736 64 0 0 37 33 0 736 64 0 0 38 0 0 736 64 0 0 38 1 0 64 32 0 0 38 2 0 288 32 0 0 38 3 0 704 64 0 0 38 4 0 480 64 0 0 38 5 0 736 64 0 0 38 6 0 736 64 0 0 38 7 0 736 64 0 0 38 8 0 736 64 0 0 38 9 0 736 64 0 0 38 10 0 736 64 0 0 38 11 0 736 64 0 0 38 12 0 736 64 0 0 38 13 0 736 64 0 0 38 14 0 736 64 0 0 38 15 0 736 64 0 0 38 16 0 736 64 0 0 38 17 0 736 64 0 0 38 18 0 736 64 0 0 38 19 0 736 64 0 0 38 20 0 736 64 0 0 38 21 0 736 64 0 0 38 22 0 736 64 0 0 38 23 0 736 64 0 0 38 24 0 736 64 0 0 38 25 0 736 64 0 0 38 26 0 736 64 0 0 38 27 0 736 64 0 0 38 28 0 736 64 0 0 38 29 0 736 64 0 0 38 30 0 736 64 0 0 38 31 0 736 64 0 0 38 32 0 736 64 0 0 38 33 0 736 64 0 0 39 0 0 704 64 0 0 39 1 0 736 64 0 0 39 2 0 288 32 0 0 39 3 0 704 64 0 0 39 4 0 512 64 0 0 39 5 0 288 64 0 0 39 6 0 288 64 0 0 39 7 0 288 64 0 0 39 8 0 288 64 0 0 39 9 0 288 64 0 0 39 10 0 512 32 0 0 39 11 0 288 64 0 0 39 12 0 288 64 0 0 39 13 0 480 64 0 0 39 14 0 544 64 0 0 39 15 0 608 0 0 0 39 16 0 576 64 0 0 39 17 0 576 64 0 0 39 18 0 576 64 1 1 40 0 0 736 64 0 0 40 1 0 480 64 0 0 40 2 0 512 64 0 0 40 3 0 512 64 0 0 40 4 0 512 64 0 0 40 5 0 288 64 0 0 40 6 0 288 64 0 0 40 7 0 288 64 0 0 40 8 0 288 64 0 0 40 9 0 512 32 0 0 40 10 0 288 64 0 0 40 11 0 288 64 0 0 40 12 0 288 64 0 0 40 13 0 288 64 0 0 40 14 0 608 0 0 0 40 15 0 544 128 0 0 40 16 0 448 0 1 0 40 17 0 448 0 1 0 40 18 0 448 0 1 1 40 19 0 448 0 1 0 40 20 0 448 0 1 0 41 0 0 736 64 0 0 41 1 0 512 64 0 0 41 2 0 288 32 0 0 41 3 0 512 96 0 0 41 4 0 512 96 0 0 41 5 0 288 64 0 0 41 6 0 768 64 0 0 41 7 0 288 64 0 0 41 8 0 480 64 0 0 41 9 0 288 64 0 0 41 10 0 288 64 0 0 41 11 0 480 64 0 0 41 12 0 288 64 0 0 41 13 0 288 64 0 0 41 14 0 512 128 0 0 41 15 0 448 0 1 0 41 16 0 448 0 1 0 41 17 0 448 0 1 0 41 18 0 448 0 1 0 41 19 0 448 0 1 0 41 20 0 448 0 1 0 42 0 0 736 64 0 0 42 1 0 512 64 0 0 42 2 0 288 32 0 0 42 3 0 512 64 0 0 42 4 0 480 64 0 0 42 5 0 288 64 0 0 42 6 0 288 64 0 0 42 7 0 768 64 0 0 42 8 0 288 64 0 0 42 9 0 768 64 0 0 42 10 0 512 32 0 0 42 11 0 288 64 0 0 42 12 0 288 64 0 0 42 13 0 544 96 0 0 42 14 0 544 128 0 0 42 15 0 448 0 1 0 42 16 0 448 0 1 0 42 17 0 448 0 1 0 42 18 0 448 0 1 0 42 19 0 448 0 1 0 42 20 0 448 0 1 0 43 0 0 736 64 0 0 43 1 0 288 32 0 0 43 2 0 512 64 0 0 43 3 0 512 96 0 0 43 4 0 512 64 0 0 43 5 0 288 64 0 0 43 6 0 288 64 0 0 43 7 0 288 64 0 0 43 8 0 768 64 0 0 43 9 0 480 64 0 0 43 10 0 480 64 0 0 43 11 0 288 64 0 0 43 12 0 288 64 0 0 43 13 0 512 128 0 0 43 14 0 448 0 1 0 43 15 0 448 0 1 0 43 16 0 448 0 1 0 43 17 0 448 0 1 0 43 18 0 448 0 1 0 43 19 0 448 0 1 0 43 20 0 448 0 1 0 44 0 0 736 64 0 0 44 1 0 512 64 0 0 44 2 0 736 96 0 0 44 3 0 512 96 0 0 44 4 0 512 64 0 0 44 5 0 288 64 0 0 44 6 0 288 64 0 0 44 7 0 288 64 0 0 44 8 0 288 64 0 0 44 9 0 480 64 0 0 44 10 0 288 64 0 0 44 11 0 288 64 0 0 44 12 0 288 64 0 0 44 13 0 512 128 0 0 44 14 0 448 0 1 0 44 15 0 448 0 1 0 44 16 0 448 0 1 0 44 17 0 448 0 1 0 44 18 0 448 0 1 0 44 19 0 448 0 1 0 44 20 0 448 0 1 0 45 0 0 736 64 0 0 45 1 0 512 64 0 0 45 2 0 736 96 0 0 45 3 0 512 64 0 0 45 4 0 512 96 0 0 45 5 0 288 64 0 0 45 6 0 288 64 0 0 45 7 0 288 64 0 0 45 8 0 480 64 0 0 45 9 0 288 64 0 0 45 10 0 288 64 0 0 45 11 0 288 64 0 0 45 12 0 544 96 0 0 45 13 0 544 128 0 0 45 14 0 448 0 1 0 45 15 0 448 0 1 0 45 16 0 448 0 1 0 45 17 0 448 0 1 0 45 18 0 448 0 1 0 45 19 0 448 0 1 0 45 20 0 448 0 1 0 46 0 0 736 64 0 0 46 1 0 288 32 0 0 46 2 0 512 64 0 0 46 3 0 736 96 0 0 46 4 0 512 64 0 0 46 5 0 288 64 0 0 46 6 0 288 64 0 0 46 7 0 288 64 0 0 46 8 0 288 64 0 0 46 9 0 288 64 0 0 46 10 0 288 64 0 0 46 11 0 288 64 0 0 46 12 0 512 128 0 0 46 13 0 448 0 1 0 46 14 0 448 0 1 0 46 15 0 448 0 1 0 46 16 0 448 0 1 0 46 17 0 448 0 1 0 46 18 0 448 0 1 0 46 19 0 448 0 1 0 46 20 0 448 0 1 0 47 0 0 736 64 0 0 47 1 0 736 96 0 0 47 2 0 288 32 0 0 47 3 0 736 96 0 0 47 4 0 480 64 0 0 47 5 0 288 64 0 0 47 6 0 288 64 0 0 47 7 0 288 64 0 0 47 8 0 288 64 0 0 47 9 0 288 64 0 0 47 10 0 288 64 0 0 47 11 0 480 64 0 0 47 12 0 512 128 0 0 47 13 0 448 0 1 0 47 14 0 448 0 1 0 47 15 0 448 0 1 0 47 16 0 448 0 1 0 47 17 0 448 0 1 0 47 18 0 448 0 1 0 47 19 0 448 0 1 0 47 20 0 448 0 1 0 48 0 0 736 64 0 0 48 1 0 512 64 0 0 48 2 0 512 64 0 0 48 3 0 512 64 0 0 48 4 0 288 32 0 0 48 5 0 288 64 0 0 48 6 0 288 64 0 0 48 7 0 64 96 0 0 48 8 0 288 64 0 0 48 9 0 288 64 0 0 48 10 0 288 64 0 0 48 11 0 288 64 0 0 48 12 0 512 128 0 0 48 13 0 448 0 1 0 48 14 0 448 0 1 0 48 15 0 448 0 1 0 48 16 0 448 0 1 0 48 17 0 448 0 1 0 48 18 0 448 0 1 0 48 19 0 448 0 1 0 48 20 0 448 0 1 0 49 0 0 736 64 0 0 49 1 0 736 96 0 0 49 2 0 480 64 0 0 49 3 0 704 64 0 0 49 4 0 512 64 0 0 49 5 0 288 64 0 0 49 6 0 288 64 0 0 49 7 0 288 64 0 0 49 8 0 288 32 0 0 49 9 0 64 96 0 0 49 10 0 288 64 0 0 49 11 0 288 64 0 0 49 12 0 640 0 0 0 49 13 0 672 64 0 0 49 14 0 672 64 0 0 49 15 0 672 64 0 0 49 16 0 704 128 0 0 49 17 0 448 0 1 0 49 18 0 448 0 1 0 49 19 0 448 0 1 0 49 20 0 448 0 1 0 50 0 0 736 64 0 0 50 1 0 736 96 0 0 50 2 0 512 64 0 0 50 3 0 512 64 0 0 50 4 0 704 64 0 0 50 5 0 288 64 0 0 50 6 0 64 96 0 0 50 7 0 288 64 0 0 50 8 0 288 64 0 0 50 9 0 288 64 0 0 50 10 0 288 32 0 0 50 11 0 288 64 0 0 50 12 0 64 32 0 0 50 13 0 288 64 0 0 50 14 0 768 64 0 0 50 15 0 288 64 0 0 50 16 0 736 128 0 0 50 17 0 448 0 1 0 50 18 0 448 0 1 0 50 19 0 448 0 1 0 50 20 0 448 0 1 0 51 0 0 736 64 0 0 51 1 0 736 96 0 0 51 2 0 512 64 0 0 51 3 0 736 96 0 0 51 4 0 512 64 0 0 51 5 0 288 64 0 0 51 6 0 288 64 0 0 51 7 0 704 64 0 0 51 8 0 288 64 0 0 51 9 0 768 64 0 0 51 10 0 288 64 0 0 51 11 0 704 64 0 0 51 12 0 288 64 0 0 51 13 0 768 64 0 0 51 14 0 288 64 0 0 51 15 0 288 64 0 0 51 16 0 736 128 0 0 51 17 0 448 0 1 0 51 18 0 448 0 1 0 51 19 0 448 0 1 0 51 20 0 448 0 1 0 52 0 0 736 64 0 0 52 1 0 512 64 0 0 52 2 0 736 96 0 0 52 3 0 480 64 0 0 52 4 0 512 64 0 0 52 5 0 288 64 0 0 52 6 0 288 64 0 0 52 7 0 288 64 0 0 52 8 0 704 64 0 0 52 9 0 32 64 0 0 52 10 0 288 64 0 0 52 11 0 768 64 0 0 52 12 0 32 64 0 0 52 13 0 288 64 0 0 52 14 0 704 64 0 0 52 15 0 32 64 0 0 52 16 0 736 128 0 0 52 17 0 448 0 1 0 52 18 0 448 0 1 0 52 19 0 448 0 1 0 52 20 0 448 0 1 0 53 0 0 736 64 0 0 53 1 0 64 32 0 0 53 2 0 480 64 0 0 53 3 0 512 64 0 0 53 4 0 704 64 0 0 53 5 0 288 64 0 0 53 6 0 288 64 0 0 53 7 0 288 32 0 0 53 8 0 288 64 0 0 53 9 0 288 64 0 0 53 10 0 704 64 0 0 53 11 0 288 64 0 0 53 12 0 704 64 0 0 53 13 0 480 64 0 0 53 14 0 288 64 0 0 53 15 0 288 64 0 0 53 16 0 736 128 0 0 53 17 0 448 0 1 0 53 18 0 448 0 1 0 53 19 0 448 0 1 0 53 20 0 448 0 1 0 54 0 0 736 64 0 0 54 1 0 512 64 0 0 54 2 0 512 64 0 0 54 3 0 64 32 0 0 54 4 0 704 64 0 0 54 5 0 288 64 0 0 54 6 0 288 64 0 0 54 7 0 288 64 0 0 54 8 0 288 64 0 0 54 9 0 480 64 0 0 54 10 0 288 64 0 0 54 11 0 64 32 0 0 54 12 0 64 32 0 0 54 13 0 288 64 0 0 54 14 0 288 64 0 0 54 15 0 480 64 0 0 54 16 0 736 128 0 0 54 17 0 448 0 1 0 54 18 0 448 0 1 0 54 19 0 448 0 1 0 54 20 0 448 0 1 0 55 0 0 448 0 1 0 55 1 0 800 64 0 0 55 2 0 800 64 0 0 55 3 0 800 64 0 0 55 4 0 768 32 0 0 55 5 0 512 96 0 0 55 6 0 512 96 0 0 55 7 0 736 32 0 0 55 8 0 768 96 0 0 55 9 0 800 64 0 0 55 10 0 800 64 0 0 55 11 0 800 64 0 0 55 12 0 800 64 0 0 55 13 0 800 64 0 0 55 14 0 800 64 0 0 55 15 0 800 64 0 0 55 16 0 768 128 0 0 55 17 0 448 0 1 0 55 18 0 448 0 1 0 55 19 0 448 0 1 0 55 20 0 448 0 1 0 56 0 0 448 0 1 0 56 1 0 448 0 1 0 56 2 0 448 0 1 0 56 3 0 448 0 1 0 56 4 0 768 0 0 0 56 5 0 768 32 0 0 56 6 0 512 64 0 0 56 7 0 512 64 0 0 56 8 0 736 128 0 0 56 9 0 448 0 1 0 56 10 0 448 0 1 0 56 11 0 448 0 1 0 56 12 0 448 0 1 0 56 13 0 448 0 1 0 56 14 0 448 0 1 0 56 15 0 448 0 1 0 56 16 0 448 0 1 0 56 17 0 448 0 1 0 56 18 0 448 0 1 0 56 19 0 448 0 1 0 56 20 0 448 0 1 0 57 0 0 448 0 1 0 57 1 0 448 0 1 0 57 2 0 448 0 1 0 57 3 0 448 0 1 0 57 4 0 448 0 1 0 57 5 0 736 0 0 0 57 6 0 512 64 0 0 57 7 0 736 96 0 0 57 8 0 736 128 0 0 57 9 0 448 0 1 0 57 10 0 448 0 1 0 57 11 0 448 0 1 0 57 12 0 448 0 1 0 57 13 0 448 0 1 0 57 14 0 448 0 1 0 57 15 0 448 0 1 0 57 16 0 448 0 1 0 57 17 0 448 0 1 0 57 18 0 448 0 1 0 57 19 0 448 0 1 0 57 20 0 448 0 1 0 58 0 0 448 0 1 0 58 1 0 448 0 1 0 58 2 0 448 0 1 0 58 3 0 448 0 1 0 58 4 0 448 0 1 0 58 5 0 736 0 0 0 58 6 0 512 96 0 0 58 7 0 512 64 0 0 58 8 0 736 128 0 0 58 9 0 448 0 1 0 58 10 0 448 0 1 0 58 11 0 448 0 1 0 58 12 0 448 0 1 0 58 13 0 448 0 1 0 58 14 0 448 0 1 0 58 15 0 448 0 1 0 58 16 0 448 0 1 0 58 17 0 448 0 1 0 58 18 0 448 0 1 0 58 19 0 448 0 1 0 58 20 0 448 0 1 0 59 0 0 448 0 1 0 59 1 0 448 0 1 0 59 2 0 448 0 1 0 59 3 0 448 0 1 0 59 4 0 448 0 1 0 59 5 0 736 0 0 0 59 6 0 736 32 0 0 59 7 0 736 32 0 0 59 8 0 736 128 0 0 59 9 0 448 0 1 0 59 10 0 448 0 1 0 59 11 0 448 0 1 0 59 12 0 448 0 1 0 59 13 0 448 0 1 0 59 14 0 448 0 1 0 59 15 0 448 0 1 0 59 16 0 448 0 1 0 59 17 0 448 0 1 0 59 18 0 448 0 1 0 59 19 0 448 0 1 0 59 20 0 448 0 1 0 60 0 0 448 0 1 0 60 1 0 448 0 1 0 60 2 0 448 0 1 0 60 3 0 448 0 1 0 60 4 0 448 0 1 0 60 5 0 736 0 0 0 60 6 0 736 96 0 0 60 7 0 512 64 0 0 60 8 0 736 128 0 0 60 9 0 448 0 1 0 60 10 0 448 0 1 0 60 11 0 448 0 1 0 60 12 0 448 0 1 0 60 13 0 448 0 1 0 60 14 0 448 0 1 0 60 15 0 448 0 1 0 60 16 0 448 0 1 0 60 17 0 448 0 1 0 60 18 0 448 0 1 0 60 19 0 448 0 1 0 60 20 0 448 0 1 0 61 0 0 448 0 1 0 61 1 0 448 0 1 0 61 2 0 448 0 1 0 61 3 0 448 0 1 0 61 4 0 448 0 1 0 61 5 0 768 0 0 0 61 6 0 768 32 0 0 61 7 0 736 32 0 0 61 8 0 736 128 0 0 61 9 0 448 0 1 0 61 10 0 448 0 1 0 61 11 0 448 0 1 0 61 12 0 448 0 1 0 61 13 0 448 0 1 0 61 14 0 448 0 1 0 61 15 0 448 0 1 0 61 16 0 448 0 1 0 61 17 0 448 0 1 0 61 18 0 448 0 1 0 61 19 0 448 0 1 0 61 20 0 448 0 1 0 62 0 0 448 0 1 0 62 1 0 448 0 1 0 62 2 0 448 0 1 0 62 3 0 448 0 1 0 62 4 0 448 0 1 0 62 5 0 448 0 1 0 62 6 0 800 32 0 0 62 7 0 800 64 0 0 62 8 0 768 128 0 0 85 0 0 736 64 0 0 86 0 0 736 64 0 0 87 0 0 736 64 0 0 88 0 0 736 64 0 0 89 0 0 736 64 0 0 90 0 0 736 64 0 0 91 0 0 736 64 0 0 92 0 0 736 64 0 0 93 0 0 736 64 0 0 94 0 0 736 64 0 0 95 0 0 736 64 0 0 96 0 0 736 64 0 0 97 0 0 736 64 0 0 98 0 0 736 64 0 0 99 0 0 736 64 0 0 100 0 0 736 64 0 0 101 0 0 736 64 0 0 102 0 0 736 64 0 0 103 0 0 736 64 0 0 104 0 0 736 64 0 0 105 0 0 736 64 0 0 106 0 0 736 64 0 0 107 0 0 736 64 0 0 108 0 0 736 64 0 0 109 0 0 736 64 0 0 110 0 0 736 64 0 0 111 0 0 736 64 0 0 112 0 0 736 64 0 0 113 0 0 736 64 0 0 114 0 0 736 64 0 0 115 0 0 736 64 0 0 116 0 0 736 64 0 0 117 0 0 736 64 0 0 118 0 0 736 64 0 0 119 0 0 736 64 0 0 120 0 0 736 64 0 0 121 0 0 736 64 0 0 122 0 0 736 64 0 0 123 0 0 736 64 0 0 124 0 0 736 64 0 0 125 0 0 736 64 0 0 126 0 0 736 64 0 0 127 0 0 736 64 0 0 128 0 0 736 64 0 0 129 0 0 736 64 0 0 130 0 0 736 64 0 0 131 0 0 736 64 0 0 132 0 0 736 64 0 0 133 0 0 736 64 0 0 134 0 0 736 64 0 0 135 0 0 736 64 0 0 136 0 0 736 64 0 0 137 0 0 736 64 0 0 138 0 0 736 64 0 0 139 0 0 736 64 0 0 140 0 0 736 64 0 0 141 0 0 736 64 0 0 142 0 0 736 64 0 0 143 0 0 736 64 0 0 144 0 0 736 64 0 0 145 0 0 736 64 0 0 146 0 0 736 64 0 0 147 0 0 736 64 0 0 148 0 0 736 64 0 0 149 0 0 736 64 0 0 