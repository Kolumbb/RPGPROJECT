150 50
32
1
0 0 0 32 32 0 0 1 0 0 32 32 0 0 5 7 0 64 0 0 0 6 7 0 64 0 0 0 6 8 0 288 224 0 0 6 9 0 288 224 0 0 6 10 0 288 224 0 0 6 11 0 288 224 0 0 6 12 0 288 224 0 0 6 13 0 288 224 0 0 6 14 0 288 224 0 0 6 15 0 288 224 0 0 7 5 0 0 0 1 0 7 6 0 32 32 1 0 7 7 0 288 0 0 0 7 8 0 288 224 0 0 7 16 0 288 224 0 0 7 17 0 288 224 0 0 8 5 0 0 0 1 0 8 6 0 32 32 1 0 8 7 0 64 0 0 0 8 8 0 288 224 0 0 8 17 0 288 224 0 0 8 18 0 288 224 0 0 9 5 0 0 0 1 0 9 6 0 32 32 1 0 9 7 0 64 0 0 0 9 8 0 288 224 0 0 9 18 0 288 224 0 0 10 4 0 0 0 1 0 10 5 0 0 0 0 0 10 6 0 32 0 0 0 10 7 0 32 32 0 0 10 8 0 288 224 0 0 10 18 0 288 224 0 0 11 4 0 0 0 1 0 11 5 0 0 0 0 0 11 6 0 288 0 0 0 11 7 0 288 224 0 0 11 8 0 288 224 0 0 11 18 0 288 224 0 0 12 4 0 0 0 1 0 12 5 0 0 0 0 0 12 6 0 288 0 0 0 12 7 0 288 224 0 0 12 18 0 288 224 0 0 13 4 0 0 0 1 0 13 5 0 0 0 0 0 13 6 0 288 0 0 0 13 7 0 288 224 0 0 13 18 0 288 224 0 0 14 4 0 0 0 1 0 14 5 0 0 0 0 0 14 6 0 288 0 0 0 14 7 0 288 224 0 0 14 18 0 288 224 0 0 15 4 0 0 0 1 0 15 5 0 0 0 0 0 15 6 0 288 0 0 0 15 7 0 288 224 0 0 15 18 0 288 224 0 0 16 4 0 0 0 1 0 16 5 0 0 0 0 0 16 6 0 288 0 0 0 16 7 0 288 224 0 0 16 8 0 288 224 0 0 16 18 0 288 224 0 0 17 4 0 0 0 1 0 17 5 0 0 0 0 0 17 6 0 320 0 0 0 17 7 0 320 32 0 0 17 8 0 288 224 0 0 17 18 0 288 224 0 0 18 5 0 0 0 1 0 18 6 0 0 0 1 0 18 7 0 288 0 0 0 18 8 0 288 224 0 0 18 18 0 288 224 0 0 19 6 0 0 0 1 0 19 7 0 288 0 0 0 19 8 0 288 224 0 0 19 18 0 288 224 0 0 20 6 0 0 0 1 0 20 7 0 288 0 0 0 20 8 0 288 224 0 0 20 12 0 32 32 0 0 20 13 0 32 32 0 0 20 17 0 288 224 0 0 20 18 0 288 224 0 0 21 6 0 0 0 1 0 21 7 0 64 0 0 0 21 8 0 288 224 0 0 21 9 0 288 224 0 0 21 15 0 288 224 0 0 21 16 0 288 224 0 0 21 17 0 288 224 0 0 22 10 0 288 224 0 0 22 11 0 288 224 0 0 22 12 0 288 224 0 0 22 13 0 288 224 0 0 22 14 0 288 224 0 0 