150 50
32
1
0 19 0 32 32 0 0 0 20 0 32 32 0 0 1 20 0 32 32 0 0 3 21 0 32 32 0 0 5 15 0 32 32 0 0 6 15 0 32 32 0 0 7 15 0 32 32 0 0 7 21 0 32 32 0 0 8 15 0 32 32 0 0 8 21 0 32 32 0 0 9 15 0 32 32 0 0 10 15 0 32 32 0 0 12 9 0 32 32 0 0 12 10 0 32 32 0 0 12 15 0 32 32 0 0 12 21 0 32 32 0 0 13 8 0 32 32 0 0 13 11 0 32 32 0 0 14 12 0 32 32 0 0 14 15 0 32 32 0 0 15 8 0 32 32 0 0 16 13 0 32 32 0 0 16 15 0 32 32 0 0 17 13 0 32 32 0 0 17 21 0 32 32 0 0 18 7 0 32 32 0 0 18 13 0 32 32 0 0 18 14 0 32 32 0 0 19 14 0 32 32 0 0 20 13 0 32 32 0 0 20 14 0 32 32 0 0 21 7 0 32 32 0 0 21 14 0 32 32 0 0 22 7 0 32 32 0 0 22 13 0 32 32 0 0 22 14 0 32 32 0 0 23 8 0 32 32 0 0 23 14 0 32 32 0 0 23 21 0 32 32 0 0 24 9 0 32 32 0 0 24 13 0 32 32 0 0 24 14 0 32 32 0 0 25 9 0 32 32 0 0 25 10 0 32 32 0 0 25 11 0 32 32 0 0 25 12 0 32 32 0 0 25 13 0 32 32 0 0 26 13 0 32 32 0 0 26 14 0 32 32 0 0 26 19 0 32 32 0 0 27 19 0 32 32 0 0 28 14 0 32 32 0 0 28 15 0 32 32 0 0 28 16 0 32 32 0 0 28 17 0 32 32 0 0 28 18 0 32 32 0 0 